module Temporizador(
	input logic PAUSE,
	input logic RESET,
	output logic [0:3] DECIMOS,
	output logic [0:3] SEGUNDOS_UNIDADE,
	output logic [0:3] SEGUNDOS_DEZENA,
	output logic [0:3] MINUTOS,
	output logic TEMPO_ACABOU
);

// PLACEHOLDER
assign DECIMOS = 0;
assign SEGUNDOS_UNIDADE = 0;
assign SEGUNDOS_DEZENA = 0;
assign MINUTOS = 0;
assign TEMPO_ACABOU = 0;

endmodule