module Comparacao (
	input logic [0:3] A,
	input logic [0:2] B,
	input logic [0:3] TENTATIVA,
	input logic START,
	input logic ENTER,
	output logic ACERTOU_SENHA_A,
	output logic ACERTOU_SENHA_B
);

endmodule