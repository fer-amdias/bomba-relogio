-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Wed Nov 19 09:24:21 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY ProjetoFinal IS 
	PORT
	(
		KEY3 :  IN  STD_LOGIC;
		KEY0 :  IN  STD_LOGIC;
		SW3 :  IN  STD_LOGIC;
		SW2 :  IN  STD_LOGIC;
		SW1 :  IN  STD_LOGIC;
		SW0 :  IN  STD_LOGIC;
		SW17 :  IN  STD_LOGIC;
		SW16 :  IN  STD_LOGIC;
		SW15 :  IN  STD_LOGIC;
		SW14 :  IN  STD_LOGIC;
		SW13 :  IN  STD_LOGIC;
		SW12 :  IN  STD_LOGIC;
		SW11 :  IN  STD_LOGIC;
		HEX0 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX1 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX2 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX3 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX4 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX5 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX6 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX7 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		LEDG :  OUT  STD_LOGIC_VECTOR(0 TO 7);
		LEDR :  OUT  STD_LOGIC_VECTOR(17 DOWNTO 0)
	);
END ProjetoFinal;

ARCHITECTURE bdf_type OF ProjetoFinal IS 

COMPONENT temporizador
	PORT(PAUSE : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 TEMPO_ACABOU : OUT STD_LOGIC;
		 DECIMOS : OUT STD_LOGIC_VECTOR(0 TO 3);
		 MINUTOS : OUT STD_LOGIC_VECTOR(0 TO 3);
		 SEGUNDOS_DEZENA : OUT STD_LOGIC_VECTOR(0 TO 3);
		 SEGUNDOS_UNIDADE : OUT STD_LOGIC_VECTOR(0 TO 3)
	);
END COMPONENT;

COMPONENT armazenamento
	PORT(SALVAR : IN STD_LOGIC;
		 SENHAS : IN STD_LOGIC_VECTOR(0 TO 6);
		 A : OUT STD_LOGIC_VECTOR(0 TO 3);
		 B : OUT STD_LOGIC_VECTOR(0 TO 2)
	);
END COMPONENT;

COMPONENT comparacao
	PORT(START : IN STD_LOGIC;
		 ENTER : IN STD_LOGIC;
		 A : IN STD_LOGIC_VECTOR(0 TO 3);
		 B : IN STD_LOGIC_VECTOR(0 TO 2);
		 TENTATIVA : IN STD_LOGIC_VECTOR(0 TO 3);
		 ACERTOU_SENHA_A : OUT STD_LOGIC;
		 ACERTOU_SENHA_B : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT circuitoativo
	PORT(START : IN STD_LOGIC;
		 ACERTOU_SENHA_B : IN STD_LOGIC;
		 ENABLE : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT menormaiordecoder7
	PORT(MENOR_OU_MAIOR : IN STD_LOGIC;
		 OUT : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT decoder7
	PORT(In : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Out : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT explosao
	PORT(TEMPO_ACABOU : IN STD_LOGIC;
		 EXPLOSAO_HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 EXPLOSAO_HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 EXPLOSAO_HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 EXPLOSAO_HEX3 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 EXPLOSAO_HEX4 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 EXPLOSAO_HEX5 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 EXPLOSAO_HEX6 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 EXPLOSAO_HEX7 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 EXPLOSAO_LEDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
	);
END COMPONENT;

COMPONENT display7mux2
	PORT(selector : IN STD_LOGIC;
		 InputA : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		 InputB : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		 Output : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mostrartentativa
	PORT(ENABLE : IN STD_LOGIC;
		 ENTER : IN STD_LOGIC;
		 ACERTOU_SENHA_A : IN STD_LOGIC;
		 TENTATIVA : IN STD_LOGIC_VECTOR(0 TO 3);
		 TENTATIVA_HEX : OUT STD_LOGIC_VECTOR(0 TO 6)
	);
END COMPONENT;

COMPONENT extensaodebitsledr
	PORT(LEDR_IN : IN STD_LOGIC_VECTOR(0 TO 3);
		 LEDR_OUT : OUT STD_LOGIC_VECTOR(0 TO 17)
	);
END COMPONENT;

COMPONENT extensaodebitsledg
	PORT(LEDG_IN : IN STD_LOGIC;
		 LEDG_OUT : OUT STD_LOGIC_VECTOR(0 TO 7)
	);
END COMPONENT;

COMPONENT ledr18mux2
	PORT(selector : IN STD_LOGIC;
		 InputA : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
		 InputB : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
		 Output : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
	);
END COMPONENT;

COMPONENT dicaparidade
	PORT(ENABLE : IN STD_LOGIC;
		 A : IN STD_LOGIC_VECTOR(0 TO 3);
		 B : IN STD_LOGIC_VECTOR(0 TO 2);
		 BIT_PARIDADE : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT dicamenormaior
	PORT(ENABLE : IN STD_LOGIC;
		 ACERTOU_SENHA_A : IN STD_LOGIC;
		 A : IN STD_LOGIC_VECTOR(0 TO 3);
		 B : IN STD_LOGIC_VECTOR(0 TO 2);
		 TENTATIVA : IN STD_LOGIC_VECTOR(0 TO 3);
		 MENOR_OU_MAIOR : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT dicabitscorretos
	PORT(ENABLE : IN STD_LOGIC;
		 ACERTOU_SENHA_A : IN STD_LOGIC;
		 A : IN STD_LOGIC_VECTOR(0 TO 3);
		 B : IN STD_LOGIC_VECTOR(0 TO 2);
		 TENTATIVA : IN STD_LOGIC_VECTOR(0 TO 3);
		 LEDR : OUT STD_LOGIC_VECTOR(0 TO 3)
	);
END COMPONENT;

SIGNAL	BIT_PARIDADE_HEX :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC_VECTOR(0 TO 2);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC_VECTOR(0 TO 6);
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC_VECTOR(0 TO 17);
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(17 DOWNTO 0);

SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(0 TO 6);
SIGNAL	GDFX_TEMP_SIGNAL_1 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	GDFX_TEMP_SIGNAL_2 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	GDFX_TEMP_SIGNAL_3 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	GDFX_TEMP_SIGNAL_4 :  STD_LOGIC_VECTOR(0 TO 3);

BEGIN 

GDFX_TEMP_SIGNAL_0 <= (SW17 & SW16 & SW15 & SW14 & SW13 & SW12 & SW11);
GDFX_TEMP_SIGNAL_1 <= (SW3 & SW2 & SW1 & SW0);
GDFX_TEMP_SIGNAL_2 <= (SW3 & SW2 & SW1 & SW0);
GDFX_TEMP_SIGNAL_3 <= (SW3 & SW2 & SW1 & SW0);
GDFX_TEMP_SIGNAL_4 <= (SW3 & SW2 & SW1 & SW0);


b2v_inst : temporizador
PORT MAP(PAUSE => SYNTHESIZED_WIRE_55,
		 RESET => SYNTHESIZED_WIRE_56,
		 TEMPO_ACABOU => SYNTHESIZED_WIRE_60,
		 DECIMOS => SYNTHESIZED_WIRE_10,
		 MINUTOS => SYNTHESIZED_WIRE_13,
		 SEGUNDOS_DEZENA => SYNTHESIZED_WIRE_12,
		 SEGUNDOS_UNIDADE => SYNTHESIZED_WIRE_11);


b2v_inst1 : armazenamento
PORT MAP(SALVAR => SYNTHESIZED_WIRE_56,
		 SENHAS => GDFX_TEMP_SIGNAL_0,
		 A => SYNTHESIZED_WIRE_58,
		 B => SYNTHESIZED_WIRE_59);


b2v_inst10 : comparacao
PORT MAP(START => SYNTHESIZED_WIRE_56,
		 ENTER => SYNTHESIZED_WIRE_57,
		 A => SYNTHESIZED_WIRE_58,
		 B => SYNTHESIZED_WIRE_59,
		 TENTATIVA => GDFX_TEMP_SIGNAL_1,
		 ACERTOU_SENHA_A => SYNTHESIZED_WIRE_62,
		 ACERTOU_SENHA_B => SYNTHESIZED_WIRE_55);


b2v_inst12 : circuitoativo
PORT MAP(START => SYNTHESIZED_WIRE_56,
		 ACERTOU_SENHA_B => SYNTHESIZED_WIRE_55,
		 ENABLE => SYNTHESIZED_WIRE_61);


b2v_inst15 : menormaiordecoder7
PORT MAP(MENOR_OU_MAIOR => SYNTHESIZED_WIRE_9,
		 OUT => SYNTHESIZED_WIRE_31);


b2v_inst16 : decoder7
PORT MAP(In => BIT_PARIDADE_HEX,
		 Out => SYNTHESIZED_WIRE_37);



b2v_inst18 : decoder7
PORT MAP(In => SYNTHESIZED_WIRE_10,
		 Out => SYNTHESIZED_WIRE_25);


b2v_inst19 : decoder7
PORT MAP(In => SYNTHESIZED_WIRE_11,
		 Out => SYNTHESIZED_WIRE_16);


b2v_inst20 : decoder7
PORT MAP(In => SYNTHESIZED_WIRE_12,
		 Out => SYNTHESIZED_WIRE_19);


b2v_inst21 : decoder7
PORT MAP(In => SYNTHESIZED_WIRE_13,
		 Out => SYNTHESIZED_WIRE_22);


b2v_inst22 : explosao
PORT MAP(TEMPO_ACABOU => SYNTHESIZED_WIRE_60,
		 EXPLOSAO_HEX0 => SYNTHESIZED_WIRE_26,
		 EXPLOSAO_HEX1 => SYNTHESIZED_WIRE_17,
		 EXPLOSAO_HEX2 => SYNTHESIZED_WIRE_20,
		 EXPLOSAO_HEX3 => SYNTHESIZED_WIRE_23,
		 EXPLOSAO_HEX4 => SYNTHESIZED_WIRE_29,
		 EXPLOSAO_HEX5 => HEX5,
		 EXPLOSAO_HEX6 => SYNTHESIZED_WIRE_32,
		 EXPLOSAO_HEX7 => SYNTHESIZED_WIRE_38,
		 EXPLOSAO_LEDR => SYNTHESIZED_WIRE_43);


b2v_inst24 : display7mux2
PORT MAP(selector => SYNTHESIZED_WIRE_60,
		 InputA => SYNTHESIZED_WIRE_16,
		 InputB => SYNTHESIZED_WIRE_17,
		 Output => HEX1);


b2v_inst25 : display7mux2
PORT MAP(selector => SYNTHESIZED_WIRE_60,
		 InputA => SYNTHESIZED_WIRE_19,
		 InputB => SYNTHESIZED_WIRE_20,
		 Output => HEX2);


b2v_inst26 : display7mux2
PORT MAP(selector => SYNTHESIZED_WIRE_60,
		 InputA => SYNTHESIZED_WIRE_22,
		 InputB => SYNTHESIZED_WIRE_23,
		 Output => HEX3);


b2v_inst27 : display7mux2
PORT MAP(selector => SYNTHESIZED_WIRE_60,
		 InputA => SYNTHESIZED_WIRE_25,
		 InputB => SYNTHESIZED_WIRE_26,
		 Output => HEX0);


b2v_inst28 : display7mux2
PORT MAP(selector => SYNTHESIZED_WIRE_60,
		 InputA => SYNTHESIZED_WIRE_28,
		 InputB => SYNTHESIZED_WIRE_29,
		 Output => HEX4);


b2v_inst29 : display7mux2
PORT MAP(selector => SYNTHESIZED_WIRE_60,
		 InputA => SYNTHESIZED_WIRE_31,
		 InputB => SYNTHESIZED_WIRE_32,
		 Output => HEX6);


b2v_inst3 : mostrartentativa
PORT MAP(ENABLE => SYNTHESIZED_WIRE_61,
		 ENTER => SYNTHESIZED_WIRE_57,
		 ACERTOU_SENHA_A => SYNTHESIZED_WIRE_62,
		 TENTATIVA => GDFX_TEMP_SIGNAL_2,
		 TENTATIVA_HEX => SYNTHESIZED_WIRE_28);


b2v_inst30 : display7mux2
PORT MAP(selector => SYNTHESIZED_WIRE_60,
		 InputA => SYNTHESIZED_WIRE_37,
		 InputB => SYNTHESIZED_WIRE_38,
		 Output => HEX7);


b2v_inst31 : extensaodebitsledr
PORT MAP(LEDR_IN => SYNTHESIZED_WIRE_39,
		 LEDR_OUT => SYNTHESIZED_WIRE_42);


b2v_inst33 : extensaodebitsledg
PORT MAP(LEDG_IN => SYNTHESIZED_WIRE_55,
		 LEDG_OUT => LEDG);


b2v_inst34 : ledr18mux2
PORT MAP(selector => SYNTHESIZED_WIRE_60,
		 InputA => SYNTHESIZED_WIRE_42,
		 InputB => SYNTHESIZED_WIRE_43,
		 Output => LEDR);


b2v_inst5 : dicaparidade
PORT MAP(ENABLE => SYNTHESIZED_WIRE_61,
		 A => SYNTHESIZED_WIRE_58,
		 B => SYNTHESIZED_WIRE_59,
		 BIT_PARIDADE => BIT_PARIDADE_HEX(0));


SYNTHESIZED_WIRE_57 <= NOT(KEY3);



SYNTHESIZED_WIRE_56 <= NOT(KEY0);



b2v_inst8 : dicamenormaior
PORT MAP(ENABLE => SYNTHESIZED_WIRE_61,
		 ACERTOU_SENHA_A => SYNTHESIZED_WIRE_62,
		 A => SYNTHESIZED_WIRE_58,
		 B => SYNTHESIZED_WIRE_59,
		 TENTATIVA => GDFX_TEMP_SIGNAL_3,
		 MENOR_OU_MAIOR => SYNTHESIZED_WIRE_9);


b2v_inst9 : dicabitscorretos
PORT MAP(ENABLE => SYNTHESIZED_WIRE_61,
		 ACERTOU_SENHA_A => SYNTHESIZED_WIRE_62,
		 A => SYNTHESIZED_WIRE_58,
		 B => SYNTHESIZED_WIRE_59,
		 TENTATIVA => GDFX_TEMP_SIGNAL_4,
		 LEDR => SYNTHESIZED_WIRE_39);


BIT_PARIDADE_HEX(2) <= '0';
BIT_PARIDADE_HEX(1) <= '0';
BIT_PARIDADE_HEX(3) <= '0';
END bdf_type;