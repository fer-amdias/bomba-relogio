module Temporizador(
	input logic PAUSE,
	input logic RESET,
	output logic [0:3] DECIMOS,
	output logic [0:3] SEGUNDOS_UNIDADE,
	output logic [0:3] SEGUNDOS_DEZENA,
	output logic [0:3] MINUTOS,
	output logic TEMPO_ACABOU
);

endmodule