module Armazenamento (
	input logic [0:6] SENHAS, 
	input logic SALVAR,
	output logic [0:3] A,
	output logic [0:2] B
);

endmodule