module Explosao(
	input logic TEMPO_ACABOU,
	input logic CLOCK,
	output logic [6:0] EXPLOSAO_HEX0,
	output logic [6:0] EXPLOSAO_HEX1,
	output logic [6:0] EXPLOSAO_HEX2,
	output logic [6:0] EXPLOSAO_HEX3,
	output logic [6:0] EXPLOSAO_HEX4,
	output logic [6:0] EXPLOSAO_HEX5,
	output logic [6:0] EXPLOSAO_HEX6,
	output logic [6:0] EXPLOSAO_HEX7,
	output logic [17:0] EXPLOSAO_LEDR
);

logic [1:0] counter; //teste
logic [1:0] counter;
logic [6:0] EXPLOSAO_HEX;
logic EXPLOSAO_LEDR0;
logic EXPLOSAO_LEDR1;
logic EXPLOSAO_LEDR2;
logic EXPLOSAO_LEDR3;

always_ff @(posedge CLOCK) begin

	if (TEMPO_ACABOU) begin
		counter <= counter + 1;
		
		if (counter == 0) begin
			EXPLOSAO_HEX[1:0]   <= 0;
			EXPLOSAO_LEDR3   <= 0;
			EXPLOSAO_LEDR2   <= 0;
			EXPLOSAO_LEDR1   <= 0;
			EXPLOSAO_LEDR0   <= 1;
			EXPLOSAO_HEX[6:2]   <= 5'b11111;
		end
		else if (counter == 1) begin
			EXPLOSAO_HEX[3:2]   <= 0;
			EXPLOSAO_LEDR3   <= 0;
			EXPLOSAO_LEDR2   <= 0;
			EXPLOSAO_LEDR1   <= 1;
			EXPLOSAO_LEDR0   <= 0;
			EXPLOSAO_HEX[6:4] <= 3'b111;
			EXPLOSAO_HEX[1:0]   <= 2'b11;
		end
		else if (counter == 2) begin
			EXPLOSAO_HEX[5:4]   <= 0;
			EXPLOSAO_LEDR3   <= 0;
			EXPLOSAO_LEDR2   <= 1;
			EXPLOSAO_LEDR1   <= 0;
			EXPLOSAO_LEDR0   <= 0;
			EXPLOSAO_HEX[6] <= 1'b1;
			EXPLOSAO_HEX[3:0]   <= 4'b1111;
		end
		else if (counter == 3) begin
			EXPLOSAO_HEX[6]   <= 0;
			EXPLOSAO_LEDR3   <= 1;
			EXPLOSAO_LEDR2   <= 0;
			EXPLOSAO_LEDR1   <= 0;
			EXPLOSAO_LEDR0   <= 0;
			EXPLOSAO_HEX[5:0] <= 6'b111111;
		end
		
			EXPLOSAO_HEX0 <= EXPLOSAO_HEX;
			EXPLOSAO_HEX1 <= EXPLOSAO_HEX;
			EXPLOSAO_HEX2 <= EXPLOSAO_HEX;
			EXPLOSAO_HEX3 <= EXPLOSAO_HEX;
			EXPLOSAO_HEX4 <= EXPLOSAO_HEX;
			EXPLOSAO_HEX5 <= EXPLOSAO_HEX;
			EXPLOSAO_HEX6 <= EXPLOSAO_HEX;
			EXPLOSAO_HEX7 <= EXPLOSAO_HEX;
			EXPLOSAO_LEDR[0]   <= EXPLOSAO_LEDR0;
			EXPLOSAO_LEDR[4]   <= EXPLOSAO_LEDR0;
			EXPLOSAO_LEDR[8]   <= EXPLOSAO_LEDR0;
			EXPLOSAO_LEDR[12]  <= EXPLOSAO_LEDR0;
			EXPLOSAO_LEDR[16]  <= EXPLOSAO_LEDR0;
			EXPLOSAO_LEDR[1]   <= EXPLOSAO_LEDR1;
			EXPLOSAO_LEDR[5]   <= EXPLOSAO_LEDR1;
			EXPLOSAO_LEDR[9]   <= EXPLOSAO_LEDR1;
			EXPLOSAO_LEDR[13]  <= EXPLOSAO_LEDR1;
			EXPLOSAO_LEDR[17]  <= EXPLOSAO_LEDR1;
			EXPLOSAO_LEDR[2]   <= EXPLOSAO_LEDR2;
			EXPLOSAO_LEDR[6]   <= EXPLOSAO_LEDR2;
			EXPLOSAO_LEDR[10]  <= EXPLOSAO_LEDR2;
			EXPLOSAO_LEDR[14]  <= EXPLOSAO_LEDR2;
			EXPLOSAO_LEDR[3]   <= EXPLOSAO_LEDR3;
			EXPLOSAO_LEDR[7]   <= EXPLOSAO_LEDR3;
			EXPLOSAO_LEDR[11]  <= EXPLOSAO_LEDR3;
			EXPLOSAO_LEDR[15]  <= EXPLOSAO_LEDR3;

	end
end

endmodule
