module MostrarTentativa (
	input logic ENABLE,
	input logic ENTER,
	input logic [0:3] TENTATIVA,
	input logic ACERTOU_SENHA_A,
	output logic [0:6] TENTATIVA_HEX
);

endmodule