module DicaMenorMaior (
	input logic ENABLE,
	input logic [0:3] TENTATIVA,
	input logic [0:3] A,
	input logic [0:2] B,
	input logic ACERTOU_SENHA_A,
	output logic MENOR_OU_MAIOR
);

endmodule