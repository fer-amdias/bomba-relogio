module Explosao(
	input logic TEMPO_ACABOU,
	output logic [6:0] EXPLOSAO_HEX0,
	output logic [6:0] EXPLOSAO_HEX1,
	output logic [6:0] EXPLOSAO_HEX2,
	output logic [6:0] EXPLOSAO_HEX3,
	output logic [6:0] EXPLOSAO_HEX4,
	output logic [6:0] EXPLOSAO_HEX5,
	output logic [6:0] EXPLOSAO_HEX6,
	output logic [6:0] EXPLOSAO_HEX7,
	output logic [17:0] EXPLOSAO_LEDR
);

endmodule
